magic
tech sky130A
magscale 1 2
timestamp 1600224028
<< error_p >>
rect 1199 1099 1210 1110
rect 1295 1099 1306 1110
rect 2524 1080 2535 1091
rect 2543 1080 2554 1091
rect 1188 726 1199 737
rect 1306 726 1317 737
rect 2554 718 2560 1080
rect 3737 975 3777 1101
rect 7217 1032 7226 1036
rect 7417 1032 7428 1043
rect 7463 1032 7474 1043
rect 6238 985 6249 996
rect 6284 985 6295 996
rect 5433 972 5444 983
rect 5479 972 5490 983
rect 3737 937 3748 948
rect 3766 937 3777 948
rect 4433 938 4444 949
rect 4479 938 4490 949
rect 3726 901 3737 912
rect 3777 901 3788 912
rect 3737 737 3777 848
rect 5433 833 5445 972
rect 7271 872 7280 1032
rect 8289 1019 8300 1030
rect 8335 1019 8346 1030
rect 7406 868 7417 879
rect 7474 868 7485 879
rect 8278 855 8289 866
rect 8346 855 8357 866
rect 6227 821 6238 832
rect 6295 821 6306 832
rect 5422 808 5433 819
rect 5490 808 5501 819
rect 4422 774 4433 785
rect 4490 774 4501 785
rect 2513 707 2524 718
rect 2554 707 2565 718
<< nwell >>
rect 879 452 1792 1358
rect 2127 433 3040 1339
rect 3341 1032 5972 1317
rect 6674 1032 7747 1317
rect 3341 411 7747 1032
rect 8102 411 9058 1317
<< varactor >>
rect 1199 726 1306 1099
rect 2524 707 2554 1080
rect 3737 901 3777 937
rect 4433 774 4490 938
rect 5433 808 5490 972
rect 6238 821 6295 985
rect 7417 868 7474 1032
rect 8289 855 8346 1019
<< pdiff >>
rect 8500 843 8621 1029
<< nsubdiff >>
rect 1047 726 1199 1099
rect 1306 726 1450 1099
rect 1653 964 1749 989
rect 1653 844 1749 869
rect 2372 707 2524 1080
rect 2554 707 2698 1080
rect 2901 945 2997 970
rect 3585 901 3737 937
rect 3777 901 3921 937
rect 4115 923 4211 948
rect 7130 992 7226 1036
rect 2901 825 2997 850
rect 4115 803 4211 828
rect 4376 774 4433 938
rect 4490 774 4572 938
rect 5299 928 5433 972
rect 5395 833 5433 928
rect 5299 808 5433 833
rect 5490 808 5572 972
rect 6181 821 6238 985
rect 6295 821 6377 985
rect 7130 872 7226 897
rect 7271 988 7417 1032
rect 7367 893 7417 988
rect 7271 868 7417 893
rect 7474 868 7556 1032
rect 8223 855 8289 1019
rect 8346 855 8428 1019
rect 8808 967 8904 1011
rect 8808 847 8904 872
<< nsubdiffcont >>
rect 1653 869 1749 964
rect 2901 850 2997 945
rect 4115 828 4211 923
rect 5299 833 5395 928
rect 7130 897 7226 992
rect 7271 893 7367 988
rect 8808 872 8904 967
<< poly >>
rect 1199 1099 1306 1259
rect 2524 1080 2554 1240
rect 1199 566 1306 726
rect 3737 937 3777 975
rect 4433 938 4490 999
rect 5433 972 5490 1033
rect 6238 985 6295 1046
rect 7417 1032 7474 1093
rect 3737 848 3777 901
rect 8289 1019 8346 1080
rect 7417 825 7474 868
rect 4433 731 4490 774
rect 5433 765 5490 808
rect 6238 778 6295 821
rect 8289 812 8346 855
rect 2524 547 2554 707
<< locali >>
rect 7130 992 7226 1036
rect 1653 964 1749 989
rect 1653 844 1749 869
rect 2901 945 2997 970
rect 2901 825 2997 850
rect 4115 923 4211 948
rect 4115 803 4211 828
rect 5299 928 5395 972
rect 7130 872 7226 897
rect 7271 988 7367 1032
rect 7271 868 7367 893
rect 8808 967 8904 1011
rect 8808 847 8904 872
rect 5299 808 5395 833
<< labels >>
flabel comment s 1390 1492 1396 1492 0 FreeSans 560 0 0 0 Incorrect:_flags_poly.5
flabel comment s 2547 304 2547 304 0 FreeSans 560 0 0 0 varac.1
flabel comment s 292 2248 292 2248 0 FreeSans 800 0 0 0 Varactor_(varac)
flabel comment s 3761 282 3761 282 0 FreeSans 560 0 0 0 varac.2
flabel comment s 1626 2208 1626 2208 0 FreeSans 560 0 0 0 Use_cif_see_NPLUS
flabel comment s 3202 2218 3202 2218 0 FreeSans 560 0 0 0 Use_cif_see_HVTP
flabel comment s 4483 311 4483 311 0 FreeSans 560 0 0 0 varac.3
flabel comment s 5329 297 5329 297 0 FreeSans 560 0 0 0 varac.4
flabel comment s 6299 283 6299 283 0 FreeSans 560 0 0 0 varac.5
flabel comment s 7243 309 7243 309 0 FreeSans 560 0 0 0 varac.6
flabel comment s 8369 315 8369 315 0 FreeSans 560 0 0 0 varac.7
flabel comment s 6270 607 6270 607 0 FreeSans 560 0 0 0 (not_implemented)
flabel comment s 8576 627 8576 627 0 FreeSans 560 0 0 0 (not_implemented)
flabel comment s -23 575 -17 575 0 FreeSans 560 0 0 0 Correct_by_design
flabel comment s -15 1143 -9 1143 0 FreeSans 560 0 0 0 Not_Implemented
flabel comment s -112 1013 -112 1013 0 FreeSans 560 0 0 0 varac.8
<< end >>
