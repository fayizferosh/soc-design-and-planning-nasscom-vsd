magic
tech sky130A
magscale 1 2
timestamp 1599840656
<< error_p >>
rect 1930 2443 2032 3111
rect 3084 2401 3089 3148
rect 3144 2404 3149 3151
rect 3189 2439 3209 3107
rect 6007 2389 6021 3113
rect 6035 2417 6049 3085
rect 1903 1547 1904 1548
rect 2275 1547 2276 1548
rect 1902 1546 2277 1547
rect 1903 1535 2276 1546
rect 1903 947 1922 1535
rect 2265 947 2276 1535
rect 2912 1486 2913 1487
rect 3196 1486 3197 1487
rect 2911 1485 2912 1486
rect 3197 1485 3198 1486
rect 3223 1306 3268 1486
rect 3477 1192 3522 1306
rect 4784 1035 4785 1036
rect 4783 1034 4784 1035
rect 2911 968 2912 969
rect 3197 968 3198 969
rect 2912 967 2913 968
rect 3196 967 3197 968
rect 1903 932 2276 947
rect 1902 931 2277 932
rect 1903 930 1904 931
rect 2275 930 2276 931
<< metal1 >>
rect 6046 989 6060 1050
rect 6121 989 6157 1050
<< via1 >>
rect 6060 989 6121 1050
<< metal2 >>
rect 3462 1192 3477 1306
rect 3574 1192 3618 1306
rect 6060 1050 6121 1111
rect 6060 923 6121 989
<< via2 >>
rect 3477 1192 3574 1306
<< metal3 >>
rect 1587 2408 1978 3155
rect 2573 2401 3089 3148
rect 3144 2404 3660 3151
rect 4299 2367 4815 3114
rect 4876 2370 5432 3117
rect 6021 2382 6506 3129
rect 1837 872 2353 1619
rect 2800 852 3316 1599
rect 3473 1306 3579 1342
rect 3473 1192 3477 1306
rect 3574 1192 3579 1306
rect 3473 1145 3579 1192
rect 4316 817 4999 1564
rect 5533 772 6049 1519
<< mimcap >>
rect 1632 2443 1930 3111
rect 2618 2436 3041 3104
rect 3189 2439 3612 3107
rect 4344 2402 4767 3070
rect 4973 2405 5384 3073
rect 6035 2417 6458 3085
rect 1882 1547 2305 1575
rect 1882 931 1903 1547
rect 2276 931 2305 1547
rect 1882 907 2305 931
rect 2845 1486 3268 1555
rect 2845 968 2912 1486
rect 3197 968 3268 1486
rect 2845 887 3268 968
rect 4361 1035 4962 1465
rect 4361 852 4784 1035
rect 5578 807 6001 1475
<< mimcapcontact >>
rect 1903 931 2276 1547
rect 2912 968 3197 1486
<< labels >>
flabel comment s 574 2516 580 2516 0 FreeSans 560 0 0 0 Correct_by_design
flabel comment s 510 2232 510 2232 0 FreeSans 560 0 0 0 mcon.3
flabel comment s 536 2059 536 2059 0 FreeSans 560 0 0 0 mcon.4
flabel comment s 393 3188 393 3188 0 FreeSans 800 0 0 0 Capm
flabel comment s 1725 2285 1725 2285 0 FreeSans 560 0 0 0 capm.1
flabel comment s 3141 2249 3141 2249 0 FreeSans 560 0 0 0 capm.2a
flabel comment s 4938 2245 4938 2245 0 FreeSans 560 0 0 0 capm.2b
flabel comment s 4836 3232 4836 3232 0 FreeSans 560 0 0 0 Incorrect
flabel comment s 6227 2303 6227 2303 0 FreeSans 560 0 0 0 capm.3
flabel comment s 520 1215 520 1215 0 FreeSans 560 0 0 0 Not required?
flabel comment s 587 1019 587 1019 0 FreeSans 560 0 0 0 capm.10
flabel comment s 596 1605 596 1605 0 FreeSans 560 0 0 0 capm.6
flabel comment s 540 1770 540 1770 0 FreeSans 560 0 0 0 Not implemented
flabel comment s 592 1439 592 1439 0 FreeSans 560 0 0 0 capm.12
flabel comment s 2088 798 2088 798 0 FreeSans 560 0 0 0 capm.4
flabel comment s 3340 792 3340 792 0 FreeSans 560 0 0 0 capm.5
flabel comment s 4737 737 4737 737 0 FreeSans 560 0 0 0 capm.7
flabel comment s 5876 693 5876 693 0 FreeSans 560 0 0 0 capm.8
flabel comment s 5779 1644 5779 1644 0 FreeSans 560 0 0 0 Incorrect
flabel comment s 5868 571 5868 571 0 FreeSans 560 0 0 0 capm.11
<< end >>
