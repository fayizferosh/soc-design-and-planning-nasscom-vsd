magic
tech sky130A
magscale 1 2
timestamp 1600224078
<< error_p >>
rect 2638 1968 2676 1972
rect 1288 1530 1298 1948
rect 1502 1530 1516 1948
rect 2667 1828 2676 1968
rect 2692 1828 2730 1968
rect 2700 1602 2734 1746
rect 3294 1624 3314 1738
rect 4228 1589 4313 1614
rect 4760 1591 4771 1616
rect 4228 1554 4288 1589
rect 5184 1358 5284 1396
rect 5764 1338 5858 1354
rect 1288 828 1298 1214
rect 1502 828 1516 1214
rect 2688 1062 2718 1190
rect 4220 1105 4280 1140
rect 2688 876 2714 1004
rect 3312 978 3344 1092
rect 4220 1080 4305 1105
rect 4810 1072 4823 1097
rect 5222 766 5316 780
rect 5784 764 5872 780
rect 5186 730 5352 744
rect 5748 728 5908 744
<< nwell >>
rect 1126 744 6196 1328
<< nmos >>
rect 2100 1708 2144 1744
<< pmos >>
rect 2148 1018 2192 1054
<< ndiff >>
rect 1268 1530 1288 1948
rect 2100 1744 2144 1902
rect 2592 1828 2676 1972
rect 2100 1584 2144 1708
rect 2596 1602 2680 1746
rect 2700 1602 2784 1746
rect 3112 1624 3256 1738
rect 3564 1626 3682 1740
rect 3722 1626 3840 1740
rect 4166 1614 4288 1728
rect 4624 1616 4746 1730
rect 5184 1358 5284 1446
<< pdiff >>
rect 1268 828 1288 1214
rect 2148 1054 2192 1194
rect 2590 1054 2664 1182
rect 2688 1062 2762 1190
rect 2148 876 2192 1018
rect 2586 868 2660 996
rect 3142 978 3286 1092
rect 3600 984 3702 1098
rect 3744 984 3862 1098
rect 4172 982 4280 1080
rect 4704 978 4798 1072
rect 5222 766 5316 860
<< psubdiff >>
rect 1486 1530 1502 1948
rect 1694 1856 1834 1880
rect 2692 1824 2776 1968
rect 5538 1816 5678 1840
rect 1694 1660 1834 1684
rect 3256 1624 3294 1738
rect 3682 1626 3722 1740
rect 4288 1576 4388 1728
rect 4746 1616 4850 1730
rect 5538 1620 5678 1644
rect 4760 1582 4850 1616
rect 5764 1338 5858 1428
<< nsubdiff >>
rect 1486 828 1502 1214
rect 1718 1116 1858 1140
rect 1718 920 1858 944
rect 2688 876 2762 1004
rect 3286 978 3312 1092
rect 3702 984 3744 1098
rect 4280 982 4372 1136
rect 4810 1072 4896 1148
rect 4798 978 4896 1072
rect 5542 1140 5682 1164
rect 5542 944 5682 968
rect 5784 764 5872 858
<< psubdiffcont >>
rect 1694 1684 1834 1856
rect 5538 1644 5678 1816
<< nsubdiffcont >>
rect 1718 944 1858 1116
rect 5542 968 5682 1140
<< poly >>
rect 2052 1708 2100 1744
rect 2144 1708 2202 1744
rect 2100 1018 2148 1054
rect 2192 1018 2232 1054
<< locali >>
rect 1694 1856 1834 1880
rect 1694 1660 1834 1684
rect 5538 1816 5678 1840
rect 5538 1620 5678 1644
rect 5542 1140 5682 1164
rect 1718 1116 1858 1140
rect 5542 944 5682 968
rect 1718 920 1858 944
<< labels >>
flabel comment s 292 2248 292 2248 0 FreeSans 800 0 0 0 Diff/tap
flabel comment s 1456 434 1456 434 0 FreeSans 560 0 0 0 difftap.1
flabel comment s 2122 1426 2122 1426 0 FreeSans 560 0 0 0 Incorrect
flabel comment s 2170 474 2170 474 0 FreeSans 560 0 0 0 difftap.2
flabel comment s 2708 456 2708 456 0 FreeSans 560 0 0 0 difftap.3
flabel comment s 3234 468 3234 468 0 FreeSans 560 0 0 0 difftap.4
flabel comment s 3740 456 3740 456 0 FreeSans 560 0 0 0 difftap.5
flabel comment s 4778 466 4782 468 0 FreeSans 560 0 0 0 difftap.7
flabel comment s 4260 472 4260 472 0 FreeSans 560 0 0 0 difftap.6
flabel comment s 5256 492 5256 492 0 FreeSans 560 0 0 0 difftap.8
flabel comment s 5226 1548 5226 1548 0 FreeSans 560 0 0 0 difftap.9
flabel comment s 5812 504 5812 504 0 FreeSans 560 0 0 0 difftap.10
flabel comment s 5814 1512 5814 1512 0 FreeSans 560 0 0 0 difftap.11
flabel comment s -16 1274 -16 1274 0 FreeSans 560 0 0 0 difftap.12
flabel comment s -22 1108 -22 1108 0 FreeSans 560 0 0 0 difftap.13
flabel comment s -18 1488 -18 1488 0 FreeSans 560 0 0 0 Unimplemented
flabel comment s 3706 1474 3706 1474 0 FreeSans 560 0 0 0 Incorrect
<< end >>
